//3
module decode (input [6:0] in, output reg [12:0] out);

	always @(in)
		begin
			case(in)
			7'b??????0: //	ANY
				out = 13'b1000000001000;
			7'b00001?1: //JC
				out = 13'b0100000001000;
			7'b00000?1: //JC
				out = 13'b1000000001000;
			7'b00011?1: //JNC
				out = 13'b1000000001000;
			7'b00010?1:	//JNC
				out = 13'b0100000001000;
			7'b0010??1: //CMPM
				out = 13'b0001001000010;
			7'b0011??1: //CMPM
				out = 13'b1001001100000;
		  	7'b0100??1: //LIT
				out = 13'b0011010000010;
			7'b0101??1: //IN
				out = 13'b0011010000100;
			7'b110??1: //LD
				out = 13'b1011010100000;
			7'b0111??1: //ST
				out = 13'b1000000111000;
			7'b1000?11: //JZ
				out = 13'b0100000001000;
			7'b1000?01: //JZ
				out = 13'b1000000001000;
			7'b1001?11: //JNZ
				out = 13'b1000000001000;
			7'b1001?01: //JNZ
				out = 13'b0100000001000;
			7'b1010??1: //ADDI
				out = 13'b0011011000010;
			7'b1011??1: //ADDM
				out = 13'b1011011100000;
			7'b1100??1: //JMP
				out = 13'b0100000001000;
			7'b1101??1: //OUT
				out = 13'b0000000001001;
		  	7'b1110??1: //NANDI
				out = 13'b0011100000010;
			7'b1111??1: //NANDM
				out = 13'b1011100100000;
			endcase
	 end
endmodule
